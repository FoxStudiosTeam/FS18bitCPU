module abstract_arithmetic_logic_unit_8bit(
    
);

endmodule