`timescale 1ns/1ps

module tb_abstract_register;

    reg clk;
    reg reset;
    reg load;
    reg [7:0] data;
    wire [7:0] current;

    // ---------------------------------------------------------
    // Генерация тактового сигнала (период 10 нс)
    // ---------------------------------------------------------
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // ---------------------------------------------------------
    // Основной тест + генерация VCD
    // ---------------------------------------------------------
    initial begin
        // --- Настройка VCD-файла ---
        $dumpfile("src/components/abstract_register/abstract_register.vcd");
        $dumpvars(0, tb_abstract_register);

        $display("=== START TEST ===");

        // Начальные значения
        reset = 1;
        load  = 0;
        data  = 8'h00;

        // Удерживаем reset некоторое время
        #12;
        reset = 0;

        // -----------------------------------------------------
        // ТЕСТ 1 — загрузка 0xA5
        // -----------------------------------------------------
        #10;
        data = 8'hA5;
        load = 1;
        #10;
        load = 0;

        // -----------------------------------------------------
        // ТЕСТ 2 — загрузка 0x3C
        // -----------------------------------------------------
        #20;
        data = 8'h3C;
        load = 1;
        #10;
        load = 0;

        // -----------------------------------------------------
        // ТЕСТ 3 — повторный reset
        // -----------------------------------------------------
        #10;
        reset = 1;
        #10;
        reset = 0;

        #20;
        data = 8'hFF;
        load = 1;
        #10;
        load =0;

        #20;
        $display("=== END TEST ===");
        $finish;
    end

    // ---------------------------------------------------------
    // Мониторинг изменений
    // ---------------------------------------------------------
    always @(posedge clk) begin
        $display("T=%0t | reset=%b load=%b data=%h -> current=%h",
                 $time, reset, load, data, current);
    end

    // ---------------------------------------------------------
    // Инстанс модуля
    // ---------------------------------------------------------
    abstract_register a_reg (
        .clk(clk),
        .reset(reset),
        .data(data),
        .load(load),
        .current(current)
    );

endmodule
